module instruction_memory (
    input [63:0] PC,     
    output reg [31:0] instruction
);
reg [7:0] memory [0:1023];


initial begin
    memory[0] = 8'h03;
    memory[1] = 8'hA4;
    memory[2] = 8'hA3;
    memory[3] = 8'h00;
    memory[4] = 8'hB3;
    memory[5] = 8'h04;
    memory[6] = 8'hA4;
    memory[7] = 8'h00;
    memory[8] = 8'h03;
    memory[9] = 8'hA4;
    memory[10] = 8'hA3;
    memory[11] = 8'h00;
    memory[12] = 8'h63;
    memory[13] = 8'h03;
    memory[14] = 8'h00;
    memory[15] = 8'h00;
    // memory[16] = 8'h23;
    // memory[17] = 8'h30;
    // memory[18] = 8'h71;
    // memory[19] = 8'h00;
    // memory[20] = 8'h03;
    // memory[21] = 8'h3F;
    // memory[22] = 8'h01;
    // memory[23] = 8'h00;
    memory[24] = 8'h23;
    memory[25] = 8'h3A;
    memory[26] = 8'h95;
    memory[27] = 8'h00;
    // memory[28] = 8'h63;
    // memory[29] = 8'h09;
    // memory[30] = 8'h00;
    // memory[31] = 8'hFE;
    // memory[32] = 8'h00;
    // memory[33] = 8'h00;
    // memory[34] = 8'h00;
    // memory[35] = 8'h00;
    // memory[36] = 8'h33;
    // memory[37] = 8'h8A;
    // memory[38] = 8'h62;
    // memory[39] = 8'h40;
    // memory[40] = 8'h63;
    // memory[41] = 8'h82;
    // memory[42] = 8'h82;
    // memory[43] = 8'h00;
    // memory[44] = 8'h33;
    // memory[45] = 8'h03;
    // memory[46] = 8'hD6;
    // memory[47] = 8'h00;
    // memory[48] = 8'hB3;
    // memory[49] = 8'h04;
    // memory[50] = 8'h83; 
    // memory[51] = 8'h40;
    // memory[52] = 8'h33;
    // memory[53] = 8'hF5;
    // memory[54] = 8'h44;
    // memory[55] = 8'h00;
    // memory[56] = 8'hB3;
    // memory[57] = 8'hE1;
    // memory[58] = 8'hA4;
    // memory[59] = 8'h00;
    // memory[60] = 8'h00;
    // memory[61] = 8'h8A;
    // memory[62] = 8'h62; 
    // memory[63] = 8'h40;
    // memory[64] = 8'h40;
    // memory[65] = 8'h40;
    // memory[66] = 8'h40;
    // memory[67] = 8'h40;
    // memory[68] = 8'h40;
    // memory[69] = 8'h40;
    // memory[70] = 8'h40;
    // memory[71] = 8'h40;
    // memory[72] = 8'h40;
    // memory[73] = 8'h40;
    // memory[74] = 8'h40;
    // memory[75] = 8'h40;
    // memory[76] = 8'h40; 
    // memory[77] = 8'h40; 
    // memory[78] = 8'h40; 
    // memory[79] = 8'h40; 
    // memory[80] = 8'hB3; 
    // memory[81] = 8'h03; 
    // memory[82] = 8'h94; 
    // memory[83] = 8'h00; 
    // memory[84] = 8'h63; 
    // memory[85] = 8'h07; 
    // memory[86] = 8'h83; 
    // memory[87] = 8'hFE; 
    // memory[88] = 8'h23; 
    // memory[89] = 8'hB1; 
    // memory[90] = 8'h62; 
    // memory[91] = 8'h00; 
    // memory[92] = 8'h03; 
    // memory[93] = 8'hB4; 
    // memory[94] = 8'h22; 
    // memory[95] = 8'h00; 
    // memory[96] = 8'h63; 
    // memory[97] = 8'h0D; 
    // memory[98] = 8'h83; 
    // memory[99] = 8'hFE; 
    // memory[100] = 8'h40; 
    // memory[101] = 8'h40; 
    // memory[102] = 8'h40; 
    // memory[103] = 8'h40; 
    // memory[104] = 8'h40; 
    // memory[105] = 8'h40; 
    // memory[106] = 8'h40; 
    // memory[107] = 8'h40; 
    // memory[108] = 8'h40;    
    // memory[109] = 8'h40;    
    // memory[110] = 8'h40;    
    // memory[111] = 8'h40;    
    // memory[112] = 8'h40;    
    // memory[113] = 8'h40;    
    // memory[114] = 8'h40;    
    // memory[115] = 8'h40;    
    // memory[116] = 8'h40;    
    // memory[117] = 8'h40;        
    // memory[118] = 8'h40;        
    // memory[119] = 8'h40;        
    // memory[120] = 8'h40;        
    // memory[121] = 8'h40;        
    // memory[122] = 8'h40;        
    // memory[123] = 8'h40;        
    // memory[124] = 8'h40;        
    // memory[125] = 8'h40;        
    // memory[126] = 8'h40;        
    // memory[127] = 8'h40;        
    // memory[128] = 8'h40;        
    // memory[129] = 8'h40;        
    // memory[130] = 8'h40;        
    // memory[131] = 8'h40;        
    // memory[132] = 8'h40;        
    // memory[133] = 8'h40;        
    // memory[134] = 8'h40;        
    // memory[135] = 8'h40;        
    // memory[136] = 8'h40;
    // memory[137] = 8'h40; 
    // memory[138] = 8'h40;
    // memory[139] = 8'h40;
    // memory[140] = 8'h40;
    // memory[141] = 8'h40;
    // memory[142] = 8'h40;
    // memory[143] = 8'h40;
    // memory[144] = 8'h40;
    // memory[145] = 8'h40;
    // memory[146] = 8'h40;
    // memory[147] = 8'h40;
    // memory[148] = 8'h40;
    // memory[149] = 8'h40;
    // memory[150] = 8'h40;
    // memory[151] = 8'h40;
    // memory[152] = 8'h40;
    // memory[153] = 8'h40;
    // memory[154] = 8'h40;
    // memory[155] = 8'h40;
    // memory[156] = 8'h40;
    // memory[157] = 8'h40;
    // memory[158] = 8'h40;
    // memory[159] = 8'h40;
    // memory[160] = 8'h40;
    // memory[161] = 8'h40;
    // memory[162] = 8'h40;
    // memory[163] = 8'h40;
    // memory[164] = 8'h40;
    // memory[165] = 8'h40;
    // memory[166] = 8'h40;
    // memory[167] = 8'h40;
    // memory[168] = 8'h40;
    // memory[169] = 8'h40;
    // memory[170] = 8'h40;
    // memory[171] = 8'h40;
    // memory[172] = 8'h40;
    // memory[173] = 8'h40;
    // memory[174] = 8'h40;
    // memory[175] = 8'h40;
    // memory[176] = 8'h40;
    // memory[177] = 8'h40;
    // memory[178] = 8'h40;
    // memory[179] = 8'h40;
    // memory[180] = 8'h40;
    // memory[181] = 8'h40;
    // memory[182] = 8'h40;
    // memory[183] = 8'h40;
    // memory[184] = 8'h40;
    // memory[185] = 8'h40;
    // memory[186] = 8'h40;
    // memory[187] = 8'h40;
    // memory[188] = 8'h40;
    // memory[189] = 8'h40;
    // memory[190] = 8'h40;
    // memory[191] = 8'h40;
    // memory[192] = 8'h40;        
    // memory[193] = 8'h40;        
    // memory[194] = 8'h40;        
    // memory[195] = 8'h40;        
    // memory[196] = 8'h40;        
    // memory[197] = 8'h40;        
    // memory[198] = 8'h40;        
    // memory[199] = 8'h40;        
    // memory[200] = 8'h40;        
    // memory[201] = 8'h40;        
    // memory[202] = 8'h40;        
    // memory[203] = 8'h40;        
    // memory[204] = 8'h40;        
    // memory[205] = 8'h40;        
    // memory[206] = 8'h40;        
    // memory[207] = 8'h40;        
    // memory[208] = 8'h40;        
    // memory[209] = 8'h40;        
    // memory[210] = 8'h40;        
    // memory[211] = 8'h40;        
    // memory[212] = 8'h40;        
    // memory[213] = 8'h40;        
    // memory[214] = 8'h40;        
    // memory[215] = 8'h40;        
    // memory[216] = 8'h40;        
    // memory[217] = 8'h40;        
    // memory[218] = 8'h40;        
    // memory[219] = 8'h40;        
    // memory[220] = 8'h40;        
    // memory[221] = 8'h40;        
    // memory[222] = 8'h40;        
    // memory[223] = 8'h40;        
    // memory[224] = 8'h40;        
    // memory[225] = 8'h40;        
    // memory[226] = 8'h40;        
    // memory[227] = 8'h40;        
    // memory[228] = 8'h40;        
    // memory[229] = 8'h40;        
    // memory[230] = 8'h40;        
    // memory[231] = 8'h40;        
    // memory[232] = 8'h40;        
    // memory[233] = 8'h40;        
    // memory[234] = 8'h40;        
    // memory[235] = 8'h40;        
    // memory[236] = 8'h40;        
    // memory[237] = 8'h40;        
    // memory[238] = 8'h40;        
    // memory[239] = 8'h40;        
    // memory[240] = 8'h40;        
    // memory[241] = 8'h40;
    // memory[242] = 8'h40;
    // memory[243] = 8'h40;
    // memory[244] = 8'h40;
    // memory[245] = 8'h40;
    // memory[246] = 8'h40;
    // memory[247] = 8'h40;
    // memory[248] = 8'h40;
    // memory[249] = 8'h40;
    // memory[250] = 8'h40;
    // memory[251] = 8'h40;
    // memory[252] = 8'h40;
    // memory[253] = 8'h40;
    // memory[254] = 8'h40;        
    // memory[255] = 8'h40;        
    // memory[256] = 8'h40;        
    // memory[257] = 8'h40;        
    // memory[258] = 8'h40;        
    // memory[259] = 8'h40;        
    // memory[260] = 8'h40;        
    // memory[261] = 8'h40;        
    // memory[262] = 8'h40;        
    // memory[263] = 8'h40;        
    // memory[264] = 8'h40;        
    // memory[265] = 8'h40;        
    // memory[266] = 8'h40;        
    // memory[267] = 8'h40;        
    // memory[268] = 8'h40;        
    // memory[269] = 8'h40;        
    // memory[270] = 8'h40;        
    // memory[271] = 8'h40;        
    // memory[272] = 8'h40;        
    // memory[273] = 8'h40;        
    // memory[274] = 8'h40;        
    // memory[275] = 8'h40;        
    // memory[276] = 8'h40;        
    // memory[277] = 8'h40;        
    // memory[278] = 8'h40;        
    // memory[279] = 8'h40;        
    // memory[280] = 8'h40;        
    // memory[281] = 8'h40;        
    // memory[282] = 8'h40;        
    // memory[283] = 8'h40;        
    // memory[284] = 8'h40;        
    // memory[285] = 8'h40;        
    // memory[286] = 8'h40;        
    // memory[287] = 8'h40;        
    // memory[288] = 8'h40;        
    // memory[289] = 8'h40;        
    // memory[290] = 8'h40;        
    // memory[291] = 8'h40;        
    // memory[292] = 8'h40;        
    // memory[293] = 8'h40;        
    // memory[294] = 8'h40;        
    // memory[295] = 8'h40;        
    // memory[296] = 8'h40;        
    // memory[297] = 8'h40;        
    // memory[298] = 8'h40;        
    // memory[299] = 8'h40;        
    // memory[300] = 8'h40;        
    // memory[301] = 8'h40;        
    // memory[302] = 8'h40;        
    // memory[303] = 8'h40;        
    // memory[304] = 8'h40;        
    // memory[305] = 8'h40;        
    // memory[306] = 8'h40;        
    // memory[307] = 8'h40;        
    // memory[308] = 8'h40;
    // memory[309] = 8'h40;
    // memory[310] = 8'h40;        
    // memory[311] = 8'h40;        
    // memory[312] = 8'h40;        
    // memory[313] = 8'h40;        
    // memory[314] = 8'h40;        
    // memory[315] = 8'h40;        
    // memory[316] = 8'h40;        
    // memory[317] = 8'h40;        
    // memory[318] = 8'h40;        
    // memory[319] = 8'h40;        
    // memory[320] = 8'h40;        
    // memory[321] = 8'h40;        
    // memory[322] = 8'h40;        
    // memory[323] = 8'h40;        
    // memory[324] = 8'h40;        
    // memory[325] = 8'h40;        
    // memory[326] = 8'h40;        
    // memory[327] = 8'h40;        
    // memory[328] = 8'h40;        
    // memory[329] = 8'h40;        
    // memory[330] = 8'h40;        
    // memory[331] = 8'h40;        
    // memory[332] = 8'h40;        
    // memory[333] = 8'h40;        
    // memory[334] = 8'h40;        
    // memory[335] = 8'h40;        
    // memory[336] = 8'h40;        
    // memory[337] = 8'h40;        
    // memory[338] = 8'h40;        
    // memory[339] = 8'h40;        
    // memory[340] = 8'h40;        
    // memory[341] = 8'h40;        
    // memory[342] = 8'h40;        
    // memory[343] = 8'h40;        
    // memory[344] = 8'h40;        
    // memory[345] = 8'h40;        
    // memory[346] = 8'h40;        
    // memory[347] = 8'h40;        
    // memory[348] = 8'h40;        
    // memory[349] = 8'h40;        
    // memory[350] = 8'h40;        
    // memory[351] = 8'h40;        
    // memory[352] = 8'h40;        
    // memory[353] = 8'h40;        
    // memory[354] = 8'h40;        
    // memory[355] = 8'h40;        
    // memory[356] = 8'h40;        
    // memory[357] = 8'h40;        
    // memory[358] = 8'h40;        
    // memory[359] = 8'h40;        
    // memory[360] = 8'h40;        
    // memory[361] = 8'h40;        
    // memory[362] = 8'h40;        
    // memory[363] = 8'h40;        
    // memory[364] = 8'h40;        
    // memory[365] = 8'h40;        
    // memory[366] = 8'h40;        
    // memory[367] = 8'h40;        
    // memory[368] = 8'h40;        
    // memory[369] = 8'h40;        
    // memory[370] = 8'h40;        
    // memory[371] = 8'h40;        
    // memory[372] = 8'h40;        
    // memory[373] = 8'h40;        
    // memory[374] = 8'h40;        
    // memory[375] = 8'h40;        
    // memory[376] = 8'h40;        
    // memory[377] = 8'h40;        
    // memory[378] = 8'h40;        
    // memory[379] = 8'h40;        
    // memory[380] = 8'h40;        
    // memory[381] = 8'h40;        
    // memory[382] = 8'h40;        
    // memory[383] = 8'h40;        
    // memory[384] = 8'h40;        
    // memory[385] = 8'h40;        
    // memory[386] = 8'h40;        
    // memory[387] = 8'h40;        
    // memory[388] = 8'h40;        
    // memory[389] = 8'h40;        
    // memory[390] = 8'h40;        
    // memory[391] = 8'h40;        
    // memory[392] = 8'h40;        
    // memory[393] = 8'h40;        
    // memory[394] = 8'h40;        
    // memory[395] = 8'h40;        
    // memory[396] = 8'h40;        
    // memory[397] = 8'h40;        
    // memory[398] = 8'h40;        
    // memory[399] = 8'h40;        
    // memory[400] = 8'h40;        
    // memory[401] = 8'h40;        
    // memory[402] = 8'h40;        
    // memory[403] = 8'h40;        
    // memory[404] = 8'h40;        
    // memory[405] = 8'h40;        
    // memory[406] = 8'h40;        
    // memory[407] = 8'h40;        
    // memory[408] = 8'h40;        
    // memory[409] = 8'h40;        
    // memory[410] = 8'h40;        
    // memory[411] = 8'h40;        
    // memory[412] = 8'h40;        
    // memory[413] = 8'h40;        
    // memory[414] = 8'h40;        
    // memory[415] = 8'h40;        
    // memory[416] = 8'h40;        
    // memory[417] = 8'h40;        
    // memory[418] = 8'h40;        
    // memory[419] = 8'h40;        
    // memory[420] = 8'h40;        
    // memory[421] = 8'h40;        
    // memory[422] = 8'h40;        
    // memory[423] = 8'h40;        
    // memory[424] = 8'h40;        
    // memory[425] = 8'h40;        
    // memory[426] = 8'h40;        
    // memory[427] = 8'h40;        
    // memory[428] = 8'h40;        
    // memory[429] = 8'h40;        
    // memory[430] = 8'h40;        
    // memory[431] = 8'h40;        
    // memory[432] = 8'h40;        
    // memory[433] = 8'h40;        
    // memory[434] = 8'h40;        
    // memory[435] = 8'h40;
    
end

wire [63:0] A1,A2,A3;
wire overflow1,overflow2,overflow3;

Cla64bit add1(
    .A(PC),
    .B(64'd1),
    .Sum(A1),
    .overflow(overflow1)
);
Cla64bit add2(
    .A(PC),
    .B(64'd2),
    .Sum(A2),
    .overflow(overflow2)
);
Cla64bit add3(
    .A(PC),
    .B(64'd3),
    .Sum(A3),
    .overflow(overflow3)
);


always @(*) begin
    instruction = {memory[A3], memory[A2], memory[A1], memory[PC]};
end
endmodule